//------------------------------------------------------------------------------
//  project:       any
//
//  packages:      rndgen_pkg
//
//  description:   parametrized synthesizable random generator pkg
//                 see Xilinx xapp 052, xapp 211
//------------------------------------------------------------------------------

`ifndef RNDGEN_SVH
`define RNDGEN_SVH

`include "rndgen.pkg"

`endif // RNDGEN_SVH

